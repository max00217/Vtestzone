module main

import vsl.plot

mut plt := plot.new_plot()

plt.add_trace(
	trace_type: .histogram
	x_str: ['China', 'India', 'USA', 'Indonesia', 'Pakistan']
	y: [1411778724.0, 1379217184, 331989449, 271350000, 225200000]
)
plt.set_layout(
	title: 'Countries by population'
)
plt.show()! 